`default_nettype none
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Dump the signals to a FST file. You can view it with gtkwave or surfer.
  initial begin
    $dumpfile("tb.fst");
    $dumpvars(0, tb);
    #1;
  end

   //parameter memfile = "hello_uart_8b.hex";
   //parameter memfile = "blink.hex";
   parameter memfile = "gpio_test.hex";
   parameter memsize = 8192;
   parameter sim = 0;
   parameter debug = 0;
   parameter width = 1;
   parameter with_csr = 0;
   parameter compressed = 0;
   parameter align = compressed;

      // Comment out direct memory access - SRAM model doesn't expose mem array
    initial
    begin
        //$display("Loading RAM from %0s", firmware_file);
        $readmemh(memfile, sram_model.mem);
    end

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;

  // Replace tt_um_example with your module name:
  tt_um_ECM24_serv_soc_top    
    dut (
      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

   // Instantiate SRAM model and connect to DUT
   sram_23lc512_model# (
        .memsize(memsize)) 
      sram_model (
       .sck(uo_out[1]),
       .cs_n(uo_out[2]),
       .si(uo_out[0]),
       .so(ui_in[0])
   );



endmodule
